module not16(i, o);
   input [15:0] i;
   output [15:0] o;
   assign o = !i;
endmodule