module not1(i, o);
   input i;
   output o;
 // always
   assign  o = !i;
endmodule
